// 启动sequence，发送到 uvm 的组件（driver)
typedef uvm_sequencer # (my_transaction) my_sequencer;

// phase
